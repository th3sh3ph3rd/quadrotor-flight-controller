vlib work
vmap work work

vcom -work work -2008 ../imu/imu_pkg.vhdl
vcom -work work -2008 ../imu/imu.vhdl
vcom -work work -2008 ../control_loop/pid_types.vhdl
vcom -work work -2008 ../control_loop/control_loop_pkg.vhdl
vcom -work work -2008 ../control_loop/control_loop.vhdl
vcom -work work -2008 ../control_loop/pid.vhdl
vcom -work work -2008 ../control_loop/calc_motor_speed.vhdl

